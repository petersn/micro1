`define SRAM_ADDRESS_SIZE 16
`define SRAM_ADDRESS_IGNORED_BITS 8
`define MEMORY_WORD_SIZE 16

module memory_controller (
  input  wire                              ena,
  input  wire                              clk,
  input  wire                              rst_n,

  // Port 0
  input  wire [`SRAM_ADDRESS_SIZE - 1 : 0] mem_address0,
  input  wire [`MEMORY_WORD_SIZE - 1 : 0]  mem_write_value0,
  input  wire                              mem_write_enable0,
  output reg  [`MEMORY_WORD_SIZE - 1 : 0]  mem_read_value0,
  input  wire                              mem_request0,
  output reg                               mem_request_complete0,

  // Port 1
  input  wire [`SRAM_ADDRESS_SIZE - 1 : 0] mem_address1,
  input  wire [`MEMORY_WORD_SIZE - 1 : 0]  mem_write_value1,
  input  wire                              mem_write_enable1,
  output reg  [`MEMORY_WORD_SIZE - 1 : 0]  mem_read_value1,
  input  wire                              mem_request1,
  output reg                               mem_request_complete1,

  output reg                               sram_cs_n,
  output reg                               sram_si,
  input  wire                              sram_so
);
  reg [11:0] counter;
  reg in_flight;
  reg which_port;

  wire [`SRAM_ADDRESS_SIZE - 1 : 0] mem_address = which_port ? mem_address1 : mem_address0;
  wire [`MEMORY_WORD_SIZE - 1 : 0] mem_write_value = which_port ? mem_write_value1 : mem_write_value0;
  wire mem_write_enable = which_port ? mem_write_enable1 : mem_write_enable0;

  always @(posedge clk) begin
    if (ena) begin
      if (!rst_n) begin
        counter <= 0;
        sram_cs_n <= 1;
        in_flight <= 0;
      end else begin
        if (in_flight) begin
          sram_cs_n <= 0;
          // The first seven bits are always 0, 0, 0, 0, 0, 0, 1
          if (counter < 6) begin
            sram_si <= 0;
          end else if (counter == 6) begin
            sram_si <= 1;
          end else if (counter == 7) begin
            // Then the eighth bit is 0 if we're writing, 1 if we're reading.
            sram_si <= !mem_write_enable;
          end else if (counter < 8 + `SRAM_ADDRESS_IGNORED_BITS) begin
            sram_si <= 0;
            // sram_si <= 1;
          end else if (counter < 32) begin
            // Then the next 17 bits are the address.
            sram_si <= mem_address[`SRAM_ADDRESS_SIZE - (counter - 8 - `SRAM_ADDRESS_IGNORED_BITS) - 1];
            //sram_si <= mem_address[counter - 8 - `SRAM_ADDRESS_IGNORED_BITS];
          end else if (counter < 32 + `MEMORY_WORD_SIZE) begin
            if (mem_write_enable) begin
              // Finally we send the bits to write, if relevant.
              sram_si <= mem_write_value[counter - 32];
            end else begin
              // Otherwise we read the bits.
              // $display("Reading bit %d = %d", counter - 32, sram_so);
              if (which_port) begin
                mem_read_value1[counter - 32] <= sram_so;
              end else begin
                mem_read_value0[counter - 32] <= sram_so;
              end
            end
          end

          if (counter < 32 + `MEMORY_WORD_SIZE) begin
            counter <= counter + 1;
          end else begin
            counter <= 32 + `MEMORY_WORD_SIZE;
            if (which_port) begin
              mem_request_complete1 <= 1;
            end else begin
              mem_request_complete0 <= 1;
            end
            sram_cs_n <= 1;
            in_flight <= 0;
          end
        end else begin
          if (mem_request0 && !mem_request_complete0) begin
            counter <= 0;
            in_flight <= 1;
            which_port <= 0;
          end else if (mem_request1 && !mem_request_complete1) begin
            counter <= 0;
            in_flight <= 1;
            which_port <= 1;
          end
        end

        // Clear completion flags, if acknowledged.
        if (!mem_request0) begin
          mem_request_complete0 <= 0;
        end
        if (!mem_request1) begin
          mem_request_complete1 <= 0;
        end
      end
    end else begin
      sram_cs_n <= 1;
    end
  end
endmodule

`define CACHE_SIZE 32

// Because memory is so slow, we need a small cache in order to stand a chance.
module cache (
  input wire ena,
  input wire clk,

  // Actual memory port.
  output reg [`SRAM_ADDRESS_SIZE - 1 : 0]  mem_address,
  output reg [`MEMORY_WORD_SIZE - 1 : 0]   mem_write_value,
  output reg                               mem_write_enable,
  input  wire  [`MEMORY_WORD_SIZE - 1 : 0] mem_read_value,
  output reg                               mem_request,
  input  wire                              mem_request_complete,

  // Cache port.
  input wire [`SRAM_ADDRESS_SIZE - 1 : 0] cache_address,
  input wire [`MEMORY_WORD_SIZE - 1 : 0]  cache_write_value,
  input wire                              cache_write_enable,
  output wire [`MEMORY_WORD_SIZE - 1 : 0] cache_read_value,
  input wire                              cache_request,
  output wire                             cache_request_complete
);
  reg [15:0] cache_values [0:`CACHE_SIZE-1];
  reg [15:0] cache_addresses [0:`CACHE_SIZE-1];

  wire [5:0] hit_cache_line = (
    cache_addresses[0] == cache_address ? 0 : cache_addresses[1] == cache_address ? 1 : cache_addresses[2] == cache_address ? 2 : cache_addresses[3] == cache_address ? 3 :
    cache_addresses[4] == cache_address ? 4 : cache_addresses[5] == cache_address ? 5 : cache_addresses[6] == cache_address ? 6 : cache_addresses[7] == cache_address ? 7 :
    cache_addresses[8] == cache_address ? 8 : cache_addresses[9] == cache_address ? 9 : cache_addresses[10] == cache_address ? 10 : cache_addresses[11] == cache_address ? 11 :
    cache_addresses[12] == cache_address ? 12 : cache_addresses[13] == cache_address ? 13 : cache_addresses[14] == cache_address ? 14 : cache_addresses[15] == cache_address ? 15 :
    cache_addresses[16] == cache_address ? 16 : cache_addresses[17] == cache_address ? 17 : cache_addresses[18] == cache_address ? 18 : cache_addresses[19] == cache_address ? 19 :
    cache_addresses[20] == cache_address ? 20 : cache_addresses[21] == cache_address ? 21 : cache_addresses[22] == cache_address ? 22 : cache_addresses[23] == cache_address ? 23 :
    cache_addresses[24] == cache_address ? 24 : cache_addresses[25] == cache_address ? 25 : cache_addresses[26] == cache_address ? 26 : cache_addresses[27] == cache_address ? 27 :
    cache_addresses[28] == cache_address ? 28 : cache_addresses[29] == cache_address ? 29 : cache_addresses[30] == cache_address ? 30 : cache_addresses[31] == cache_address ? 31 : 32
  );
  // The first 4096 bytes of memory are never cached.
  wire cache_miss = hit_cache_line[5] || (cache_address < 16'h1000);

  reg [4:0] eviction_counter = 0;

  always @(posedge clk) begin
    if (ena) begin
      // Check for an incoming request to the cache.
      if (cache_request) begin
        if (cache_miss) begin
          if (cache_write_enable) begin
            // === Handle a cache miss write ===
            if (!mem_request) begin
              // Write the value to the cache.
              cache_values[eviction_counter] <= cache_write_value;
              cache_addresses[eviction_counter] <= cache_address;
              eviction_counter <= eviction_counter + 1;
              mem_request <= 1;
              mem_address <= cache_address;
              mem_write_value <= cache_write_value;
              mem_write_enable <= 1;
            end else begin
              // Pass on a response, if relevant.
              if (mem_request_complete) begin
                cache_request_complete <= 1;
              end
            end
          end else begin
            // === Handle a cache miss read ===
            if (!mem_request) begin
              // Read the value from memory.
              mem_request <= 1;
              mem_address <= cache_address;
              mem_write_enable <= 0;
            end else begin
              // Pass on a response, if relevant.
              if (mem_request_complete) begin
                cache_read_value <= mem_read_value;
                cache_request_complete <= 1;
              end
            end
          end
        end else if (!cache_request_complete) begin
          if (cache_write_enable) begin
            // === Handle a cache hit write ===
            cache_values[hit_cache_line] <= cache_write_value;
            cache_addresses[hit_cache_line] <= cache_address;
            cache_request_complete <= 1;
          end else begin
            // === Handle a cache hit read ===
            cache_read_value <= cache_values[hit_cache_line];
            cache_request_complete <= 1;
          end
        end
      end else begin
        // Otherwise, acknowledge the request.
        cache_request_complete <= 0;
      end
    end
  end
endmodule

module font_rom(
  input wire [7:0] char,
  input wire [3:0] pixel_x,
  input wire [3:0] pixel_y,
  output wire color
);
  reg [255:0] font [0:95];
  initial begin
    font[0] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    font[1] = 256'b0000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000;
    font[2] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011000000000011001100000000001100110000000000110011000;
    font[3] = 256'b0000000000000000000000000000000000000001100110000000000110011000000000011001100000000001100110000000011111111110000001111111111000000001100110000000000110011000000001111111111000000111111111100000000110011000000000011001100000000001100110000000000110011000;
    font[4] = 256'b0000000000000000000000000000000000000000011000000000000001100000000000011111111000000011111111100000011001100000000001100110000000000011111111000000000111111110000000000110011000000000011001100000011111111110000001111111110000000000011000000000000001100000;
    font[5] = 256'b0000000000000000000000000000000000000111100001100000011110000110000001111000011000000111100011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100011110000001100001111000000110000111100000011000011110;
    font[6] = 256'b0000000000000000000000000000000000000010011111000000001111111110000000111100011000000011110001100000001111100110000000100111111000000000001111000000000000111100000000000111111000000000011001100000000001100110000000000110011000000000001111100000000000011100;
    font[7] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000000011000000000000001100000;
    font[8] = 256'b0000000000000000000000000000000000000001110000000000000111100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000001111000000000000111000000;
    font[9] = 256'b0000000000000000000000000000000000000000000110000000000000111000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000001110000000000000011000;
    font[10] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011000000000011001100000000000111100000000000011110000000001111111111000000111111111100000000011110000000000001111000000000001100110000000000110011000;
    font[11] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000011000000000000001100000000000000110000000000111111111100000011111111110000000000110000000000000011000000000000001100000000000000110000000000000000000000000000000000000;
    font[12] = 256'b0000000000011000000000000011100000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    font[13] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    font[14] = 256'b0000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    font[15] = 256'b0000000000000000000000000000000000000000000001100000000000000110000000000000011000000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000001100000000000000110000000000000011000000000;
    font[16] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000011110000001100011111000000110011101100000011011100110000001111100011000000111100001100000011100000110000001100000011000000011111111100000000111111100;
    font[17] = 256'b0000000000000000000000000000000000000001111110000000000111111000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001111000000000000111100000000000011100000000000001100000;
    font[18] = 256'b0000000000000000000000000000000000000111111111100000011111111110000000000001110000000000001110000000000001110000000000001110000000000001110000000000001110000000000001110000000000000110000000000000011000000110000001100000011000000011111111100000000111111100;
    font[19] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000000000001100000000000000011111000000000001111100000000001100000000000000110000000000000011000000110000001100000011000000011111111100000000111111100;
    font[20] = 256'b0000000000000000000000000000000000000001100000000000000110000000000000011000000000000001100000000000011111111110000001111111111000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100000000000000110000000;
    font[21] = 256'b0000000000000000000000000000000000000001111111100000001111111110000001100000000000000110000000000000011000000000000001100000000000000011111111100000000111111110000000000000011000000000000001100000000000000110000000000000011000000011111111100000001111111110;
    font[22] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111110000000000000011000000000000001100000000000000110000000000000011000000001111111100000000111111100;
    font[23] = 256'b0000000000000000000000000000000000000000000000100000000000000110000000000000110000000000000111000000000000111000000000000111000000000000111000000000000111000000000000111000000000000011000000000000001100000000000000110000000000000011111111100000001111111110;
    font[24] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000001111111100000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111100;
    font[25] = 256'b0000000000000000000000000000000000000001111111100000001111111110000001100000000000000110000000000000011000000000000001100000000000000111111111000000011111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111100;
    font[26] = 256'b0000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000011110000000000001111000000000000111100000000000000000000000000000000000;
    font[27] = 256'b0000000000011000000000000011100000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000011110000000000001111000000000000111100000000000000000000000000000000000;
    font[28] = 256'b0000000000000000000000000000000000000000100000000000000011000000000000000110000000000000001100000000000000111000000000000001110000000000000011100000000000001110000000000001110000000000001110000000000000110000000000000110000000000000110000000000000010000000;
    font[29] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000000000000000000000000000000000000001111111111000000111111111100000000000000000000000000000000000000000000000000000000000000000;
    font[30] = 256'b0000000000000000000000000000000000000000000110000000000000111000000000000111000000000000111000000000000111000000000000011000000000000011000000000000001100000000000000011000000000000001110000000000000011100000000000000111000000000000001110000000000000011000;
    font[31] = 256'b0000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000000001100000000000001110000000000001110000000000001110000000000001110000000000000110000000000000011000000110000001100000011000000011111111100000000111111100;
    font[32] = 256'b0000000000000000000000000000000000000111111111000000011111111110000000000000011000000000000001100000000111000110000000111110011000000110011001100000011001100110000001111110011000000111110001100000011000000110000001100000011000000011111111100000000111111100;
    font[33] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000111111111100000011111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111100;
    font[34] = 256'b0000000000000000000000000000000000000001111111100000001111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000001111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111110;
    font[35] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000011000000110000001100000011000000011111111100000000111111100;
    font[36] = 256'b0000000000000000000000000000000000000001111111100000001111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111110;
    font[37] = 256'b0000000000000000000000000000000000000011111111100000001111111110000000000000011000000000000001100000000000000110000000000000011000000000111111100000000011111110000000000000011000000000000001100000000000000110000000000000011000000011111111100000001111111110;
    font[38] = 256'b0000000000000000000000000000000000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000111111100000000011111110000000000000011000000000000001100000000000000110000000000000011000000011111111100000001111111110;
    font[39] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000110000001100000011000000111100001100000011110000110000000000000011000000000000001100000011000000110000001100000011000000011111111100000000111111100;
    font[40] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000111111111100000011111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110;
    font[41] = 256'b0000000000000000000000000000000000000001111110000000000111111000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000001111110000000000111111000;
    font[42] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000;
    font[43] = 256'b0000000000000000000000000000000000000010000001100000001100000110000000011000011000000001110001100000000011100110000000000111111000000000001111100000000000111110000000000111011000000000111001100000000011000110000000011000011000000011000001100000001000000110;
    font[44] = 256'b0000000000000000000000000000000000000011111111100000001111111110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110;
    font[45] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100110011000000110111101100000011111111110000001111001111000000111000011100000011000000110;
    font[46] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001110000011000000111100001100000011111000110000001101110011000000110011101100000011000111110000001100001111000000110000011100000011000000110;
    font[47] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111100;
    font[48] = 256'b0000000000000000000000000000000000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000001111111100000001111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111110;
    font[49] = 256'b0000000000000000000000000000000000000110011111000000011111111110000000111100011000000011110001100000011111100110000001100110011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111100;
    font[50] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000011111111100000001111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111110;
    font[51] = 256'b0000000000000000000000000000000000000011111111000000001111111110000001100000011000000110000001100000011000000000000001100000000000000011111111000000000111111110000000000000011000000000000001100000011000000110000001100000011000000011111111100000000111111100;
    font[52] = 256'b0000000000000000000000000000000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000111111111100000011111111110;
    font[53] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110;
    font[54] = 256'b0000000000000000000000000000000000000000011000000000000011110000000000011111100000000011100111000000011100001110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110;
    font[55] = 256'b0000000000000000000000000000000000000001110111000000001111111110000001100110011000000110011001100000011001100110000001100110011000000110011001100000011001100110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110;
    font[56] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000111000011100000001110011100000000011111100000000000111100000000000011110000000000011111100000000011100111000000011100001110000001100000011000000110000001100000011000000110;
    font[57] = 256'b0000000000000000000000000000000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000011110000000000011111100000000011100111000000011100001110000001100000011000000110000001100000011000000110;
    font[58] = 256'b0000000000000000000000000000000000000011111111100000001111111110000000000000011000000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000001100000000000000111111111000000011111111100;
    font[59] = 256'b0000000000000000000000000000000000000001111000000000000111100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000001111000000000000111100000;
    font[60] = 256'b0000000000000000000000000000000000000110000000000000011000000000000001100000000000000111000000000000001110000000000000011100000000000000111000000000000001110000000000000011100000000000000111000000000000001110000000000000011000000000000001100000000000000110;
    font[61] = 256'b0000000000000000000000000000000000000000011110000000000001111000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011110000000000001111000;
    font[62] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000111000011100000001110011100000000011111100000000000111100000000000001100000;
    font[63] = 256'b0000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    font[64] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000011100000000000000111000000000000001100000;
    font[65] = 256'b0000000000000000000000000000000000000111111111000000011111111110000001100000011000000110000001100000011111111110000001111111110000000110000000000000011000000000000000111111100000000001111110000000000000000000000000000000000000000000000000000000000000000000;
    font[66] = 256'b0000000000000000000000000000000000000001111111100000001111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000000111111111000000001111111100000000000000110000000000000011000000000000001100000000000000110;
    font[67] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000000000000110000000000000011000000110000001100000011000000110000000111111111000000001111111000000000000000000000000000000000000000000000000000000000000000000;
    font[68] = 256'b0000000000000000000000000000000000000111111111000000011111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001111111111000000111111111000000011000000000000001100000000000000110000000000000011000000000;
    font[69] = 256'b0000000000000000000000000000000000000001111111000000000111111110000000000000011000000000000001100000011111111110000001111111111000000110000001100000011000000110000000111111111000000001111111000000000000000000000000000000000000000000000000000000000000000000;
    font[70] = 256'b0000000000000000000000000000000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000011111100000000001111110000000000001100000000000000110000000000011111000000000001111000000;
    font[71] = 256'b0000000111111000000000111111100000000110000000000000011000000000000001111111110000000111111111100000011000000110000001100000011000000110000001100000011000000110000001111111111000000111111111000000000000000000000000000000000000000000000000000000000000000000;
    font[72] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000000111111111000000001111111100000000000000110000000000000011000000000000001100000000000000110;
    font[73] = 256'b0000000000000000000000000000000000000001111110000000000111111000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000111100000000000011110000000000000000000000000000000000000000000011000000000000001100000;
    font[74] = 256'b0000000001111100000000001111111000000001100001100000000110000110000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011110000000000001111000000000000000000000000000000000000000000001100000000000000110000000;
    font[75] = 256'b0000000000000000000000000000000000000010000110000000001100011000000000111001100000000001111110000000000011111000000000001111100000000001110110000000001110011000000000110001100000000010000110000000000000011000000000000001100000000000000110000000000000011000;
    font[76] = 256'b0000000000000000000000000000000000000001111110000000000111111000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011110000000000001111000;
    font[77] = 256'b0000000000000000000000000000000000000110011001100000011001100110000001100110011000000110011001100000011001100110000001100110011000000110011001100000011001100110000000111111111000000001100111100000000000000000000000000000000000000000000000000000000000000000;
    font[78] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000000111111111000000001111111100000000000000000000000000000000000000000000000000000000000000000;
    font[79] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000000111111111000000001111111000000000000000000000000000000000000000000000000000000000000000000;
    font[80] = 256'b0000000000000110000000000000011000000000000001100000000000000110000000011111111000000011111111100000011000000110000001100000011000000110000001100000011000000110000000111111111000000001111111100000000000000000000000000000000000000000000000000000000000000000;
    font[81] = 256'b0000011000000000000001100000000000000110000000000000011000000000000001111111110000000111111111100000011000000110000001100000011000000110000001100000011000000110000001111111111000000111111111000000000000000000000000000000000000000000000000000000000000000000;
    font[82] = 256'b0000000000000000000000000000000000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000110000110000000011000011000000000111111100000000001111110000000000000000000000000000000000000000000000000000000000000000000;
    font[83] = 256'b0000000000000000000000000000000000000001111111100000001111111110000001100000000000000110000000000000001111111100000000011111111000000000000001100000000000000110000001111111111000000111111111000000000000000000000000000000000000000000000000000000000000000000;
    font[84] = 256'b0000000000000000000000000000000000000111110000000000011111100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000001111111100000000111111110000000000001100000000000000110000000000000011000000000000001100000;
    font[85] = 256'b0000000000000000000000000000000000000111111111000000011111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000000000000000000000000000000000000000000000000000000000000000;
    font[86] = 256'b0000000000000000000000000000000000000000011000000000000011110000000000011111100000000011100111000000011100001110000001100000011000000110000001100000011000000110000001100000011000000110000001100000000000000000000000000000000000000000000000000000000000000000;
    font[87] = 256'b0000000000000000000000000000000000000001110111000000001111111110000001100110011000000110011001100000011001100110000001100110011000000110011001100000011001100110000001100000011000000110000001100000000000000000000000000000000000000000000000000000000000000000;
    font[88] = 256'b0000000000000000000000000000000000000110000001100000011100001110000000111001110000000001111110000000000011110000000000001111000000000001111110000000001110011100000001110000111000000110000001100000000000000000000000000000000000000000000000000000000000000000;
    font[89] = 256'b0000000111111000000000111111100000000110000000000000011000000000000001111111110000000111111111100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000000000000000000000000000000000000000000000000000000000000000;
    font[90] = 256'b0000000000000000000000000000000000000111111111100000011111111110000000000001110000000000001110000000000001110000000000001110000000000001110000000000001110000000000001111111111000000111111111100000000000000000000000000000000000000000000000000000000000000000;
    font[91] = 256'b0000000000000000000000000000000000000001110000000000000111100000000000000110000000000000011000000000000001100000000000000110000000000000001110000000000000111000000000000110000000000000011000000000000001100000000000000110000000000001111000000000000111000000;
    font[92] = 256'b0000000000000000000000000000000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000;
    font[93] = 256'b0000000000000000000000000000000000000000000110000000000000111000000000000110000000000000011000000000000001100000000000000110000000000001110000000000000111100000000000000110000000000000011000000000000001100000000000000110000000000000001110000000000000011000;
    font[94] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000011111000000000011001100110000001100110011000000000001111000000000000011100;
    font[95] = 256'b0000000000000000000000000000000000000111111111100000011111111110000001111111111000000111111111100000011111111110000001111111111000000111111111100000011111111110000001111111111000000111111111100000011111111110000001111111111000000111111111100000011111111110;
  end
  assign color = ((char >= 32) && (char < 96)) ? font[char - 32][pixel_y * 16 + pixel_x] : pixel_x ^ pixel_y;
endmodule

// PMOD0 is the output for the VGA.
// PMOD1 is the input/output for the SRAM.
//   PMOD1[0]: ~CS
//   PMOD1[1]: SO
//   PMOD1[2]: SIO2
//   PMOD1[3]: SI
//   PMOD1[4]: SCK
//   PMOD1[5]: ~HOLD/SIO3

`define WORD_SIZE 16
`define REGISTER_COUNT 16

module processor(
  input  wire       ena,        // high when enabled
  input  wire       clk_100mhz, // clock
  input  wire       rst_n,       // reset negated (low to reset)

  output wire error_out, // high when an error has occurred

  // Memory port.
  output reg [`SRAM_ADDRESS_SIZE - 1 : 0]  mem_address,
  output reg [`MEMORY_WORD_SIZE - 1 : 0]   mem_write_value,
  output reg                               mem_write_enable,
  input  wire  [`MEMORY_WORD_SIZE - 1 : 0] mem_read_value,
  output reg                               mem_request,
  input  wire                              mem_request_complete
);
  // CPU state.
  reg error;
  reg [`WORD_SIZE - 1 : 0] register_file[`REGISTER_COUNT];
  reg [`SRAM_ADDRESS_SIZE - 1 : 0] instruction_pointer;
  reg [`WORD_SIZE - 1 : 0] fetched_instruction;
  reg ifetch_required;

  assign error_out = error;

  // Aliases.
  wire [3:0] regA;
  assign regA = fetched_instruction[11:8];
  wire [3:0] regB;
  assign regB = fetched_instruction[15:12];
  wire [3:0] regDest;
  assign regDest = fetched_instruction[7:4];
  wire [3:0] imm4;
  assign imm4 = fetched_instruction[15:12];
  wire [15:0] imm4SignExtended;
  assign imm4SignExtended = {{12{imm4[3]}}, imm4};
  wire [7:0] imm8;
  assign imm8 = fetched_instruction[15:8];
  wire [15:0] imm8SignExtended;
  assign imm12SignExtended = {{8{imm8[7]}}, imm8};
  wire [11:0] imm12;
  assign imm12 = fetched_instruction[15:4];
  wire [15:0] imm12SignExtended;
  assign imm12SignExtended = {{4{imm12[11]}}, imm12};

  always @(posedge clk) begin
    if (ena) begin
      if (!rst_n) begin
        error <= 0;
        instruction_pointer <= 16'h1000;
        mem_request <= 0;
        ifetch_required <= 1;
      end else if (!error) begin
        // ========== Main logic begins here ==========

        // If we don't have the instruction fetched, then fetch it.
        if (ifetch_required) begin
          mem_address <= instruction_pointer;
          mem_request <= 1;
          mem_write_enable <= 0;
          if (mem_request_complete) begin
            mem_request <= 0;
            // $display("Fetched instruction @%h %b", instruction_pointer, mem_read_value);
            fetched_instruction <= mem_read_value;
            ifetch_required <= 0;
            instruction_pointer <= instruction_pointer + 2;
          end
        end else begin
          case (fetched_instruction[3:0])
            4'b0000: begin
              // $display("HCF");
              error <= 1;
            end
            4'b0001: begin
              // Perform an unary operation.
              case (regB)
                4'b0000: begin
                  // $display("MOV r%d = r%d", regDest, regA);
                  register_file[regDest] <= register_file[regA];
                end
                4'b0001: begin
                  // $display("NOT r%d = ~r%d", regDest, regA);
                  register_file[regDest] <= ~register_file[regA];
                end
                4'b0010: begin
                  // $display("NEG r%d = -r%d", regDest, regA);
                  register_file[regDest] <= -register_file[regA];
                end
                4'b0011: begin
                  // $display("INC r%d = r%d + 1", regDest, regA);
                  register_file[regDest] <= register_file[regA] + 1;
                end
                4'b0100: begin
                  // $display("DEC r%d = r%d - 1", regDest, regA);
                  register_file[regDest] <= register_file[regA] - 1;
                end
              endcase
              ifetch_required <= 1;
            end
            4'b0010: begin
              // $display("ADD r%d = r%d + r%d", regDest, regA, regB);
              register_file[regDest] <= register_file[regA] + register_file[regB];
              ifetch_required <= 1;
            end
            4'b0011: begin
              // $display("LIT8 r%d = %d", regDest, imm8SignExtended);
              register_file[regDest] <= imm8SignExtended;
              ifetch_required <= 1;
            end
            4'b0100: begin
              // $display("LIT8H r%d = %d", regDest, imm8SignExtended);
              register_file[regDest][15:8] <= imm8;
              ifetch_required <= 1;
            end
            4'b0101: begin
              // $display("JNZ %d, r%d", $signed(imm8SignExtended), regDest);
              if (register_file[regDest] != 0) begin
                instruction_pointer <= instruction_pointer + imm8SignExtended;
              end
              ifetch_required <= 1;
            end
            4'b0110: begin
              // $display("JMP %d", $signed(imm12SignExtended));
              instruction_pointer <= instruction_pointer + imm12SignExtended;
              ifetch_required <= 1;
            end
            4'b0111: begin
              // $display("LOAD r%d = [r%d + %d]", regDest, regA, $signed(imm4SignExtended));
              mem_address <= register_file[regA] + imm4SignExtended;
              mem_request <= 1;
              mem_write_enable <= 0;
              if (mem_request_complete) begin
                // $display("Loaded %d", mem_read_value);
                mem_request <= 0;
                register_file[regDest] <= mem_read_value;
                ifetch_required <= 1;
              end
            end
            4'b1000: begin
              // $display("STORE [r%d + %d] = r%d", regA, $signed(imm4SignExtended), regB);
              mem_address <= register_file[regA] + imm4SignExtended;
              mem_write_value <= register_file[regB];
              mem_request <= 1;
              mem_write_enable <= 1;
              if (mem_request_complete) begin
                // $display("Stored");
                mem_request <= 0;
                ifetch_required <= 1;
              end
            end
            default: begin
              // $display("BADOP");
              error <= 1;
            end
          endcase
        end
      end
    end
  end
endmodule

module micro1 (
  input  wire [7:0] ui_in,      // dedicated inputs
  output wire [7:0] uo_out,     // dedicated outputs
  input  wire [7:0] uio_in,     // bidirectional input path
  output wire [7:0] uio_out,    // bidirectional output path
  output wire [7:0] uio_oe,     // bidir output enable (high=out)
  input  wire       ena,        // high when enabled
  input  wire       clk_100mhz, // clock
  input  wire       rst_n,       // reset negated (low to reset)
  output wire       led        // LED output
);
  wire vga_r = uo_out[0];
  wire vga_g = uo_out[1];
  wire vga_b = uo_out[2];
  wire vga_hs = uo_out[3];
  wire vga_vs = uo_out[4];

  reg [`SRAM_ADDRESS_SIZE - 1 : 0] video_mem_address;
  reg [`MEMORY_WORD_SIZE - 1 : 0]  video_mem_write_value;
  reg                              video_mem_write_enable;
  reg [`MEMORY_WORD_SIZE - 1 : 0]  video_mem_read_value;
  reg                              video_mem_request;
  reg                              video_mem_request_complete;

  reg [`SRAM_ADDRESS_SIZE - 1 : 0] cpu_mem_address;
  reg [`MEMORY_WORD_SIZE - 1 : 0]  cpu_mem_write_value;
  reg                              cpu_mem_write_enable;
  reg [`MEMORY_WORD_SIZE - 1 : 0]  cpu_mem_read_value;
  reg                              cpu_mem_request;
  reg                              cpu_mem_request_complete;

  reg [`SRAM_ADDRESS_SIZE - 1 : 0] cache_mem_address;
  reg [`MEMORY_WORD_SIZE - 1 : 0]  cache_mem_write_value;
  reg                              cache_mem_write_enable;
  reg [`MEMORY_WORD_SIZE - 1 : 0]  cache_mem_read_value;
  reg                              cache_mem_request;
  reg                              cache_mem_request_complete;

  // Instantiate the cache.
  cache cache_inst(
    .ena(ena),
    .clk(clk_100mhz),

    .mem_address(cpu_mem_address),
    .mem_write_value(cpu_mem_write_value),
    .mem_write_enable(cpu_mem_write_enable),
    .mem_read_value(cpu_mem_read_value),
    .mem_request(cpu_mem_request),
    .mem_request_complete(cpu_mem_request_complete),

    .cache_address(cache_mem_address),
    .cache_write_value(cache_mem_write_value),
    .cache_write_enable(cache_mem_write_enable),
    .cache_read_value(cache_mem_read_value),
    .cache_request(cache_mem_request),
    .cache_request_complete(cache_mem_request_complete)
  );

  wire error_out;
  assign led = !error_out;

  // Instantiate the main processor.
  processor processor_inst(
    .ena(ena),
    .clk_100mhz(clk_100mhz),
    .rst_n(rst_n),

    .error_out(error_out),

    .mem_address(cache_mem_address),
    .mem_write_value(cache_mem_write_value),
    .mem_write_enable(cache_mem_write_enable),
    .mem_read_value(cache_mem_read_value),
    .mem_request(cache_mem_request),
    .mem_request_complete(cache_mem_request_complete)
  );

  // Set output directions.
  assign uio_oe[0] = 1;
  assign uio_oe[1] = 0;
  assign uio_oe[2] = 1; // We're pulling up, so output.
  assign uio_oe[3] = 1;
  assign uio_oe[4] = 1;
  assign uio_oe[5] = 1; // We're pulling up, so output.
  // Assign pull-up values.
  assign uio_out[2] = 1;
  assign uio_out[5] = 1;

  reg [3:0] mem_controller_clock_divider = 0;
  always @(posedge clk_100mhz) begin
    mem_controller_clock_divider <= mem_controller_clock_divider + 1;
  end

  // Assign the serial clock.
  assign uio_out[4] = !(mem_controller_clock_divider[3] ^ mem_controller_clock_divider[2]);

  memory_controller memory_controller_inst(
    .ena(ena),
    .clk(mem_controller_clock_divider[3]),
    .rst_n(rst_n),

    .mem_address0(video_mem_address),
    .mem_write_value0(video_mem_write_value),
    .mem_write_enable0(video_mem_write_enable),
    .mem_read_value0(video_mem_read_value),
    .mem_request0(video_mem_request),
    .mem_request_complete0(video_mem_request_complete),

    .mem_address1(cpu_mem_address),
    .mem_write_value1(cpu_mem_write_value),
    .mem_write_enable1(cpu_mem_write_enable),
    .mem_read_value1(cpu_mem_read_value),
    .mem_request1(cpu_mem_request),
    .mem_request_complete1(cpu_mem_request_complete),

    .sram_cs_n(uio_out[0]),
    .sram_si(uio_out[3]),
    .sram_so(uio_in[1])
  );

  reg [23:0] ctr = 0;
  reg [15:0] scanline = 0;
  reg [31:0] lfsr = 1;

  reg [15:0] line_buffer1 [0:19];
  reg [15:0] line_buffer2 [0:19];
  reg line_flip = 0;
  reg [5:0] line_ctr = 0;
  reg [4:0] line_ptr = 0;

  reg mem_fill = 0;

  wire video_en = (scanline >= 35) && (scanline < 515) && (ctr < 2700);

  // We now figure out which character we're at.
  wire [9:0] offset_scanline = scanline - 35;
  wire [4:0] current_row = offset_scanline[8:4];
  wire [3:0] pixel_y = offset_scanline[3:0];
  // Each pixel is 4 cycles long.
  wire [6:0] current_col = ctr[12:6];
  wire [3:0] pixel_x = ctr[5:2];

  wire [15:0] current_char_pair = current_col >= 40 ? 0 : (line_flip ? line_buffer2[current_col >> 1] : line_buffer1[current_col >> 1]);
  wire [7:0] current_char = current_col[0] ? current_char_pair[7:0] : current_char_pair[15:8];

  wire color;
  font_rom font_rom_inst(
    .char(current_char),
    .pixel_x(pixel_x),
    .pixel_y(pixel_y),
    .color(color)
  );

  // We now interpret the character as a little 2x4 grid.
  // wire color = current_char[{pixel_y[3], pixel_y[2], pixel_x[3]}];
  //wire color = (current_col >= 39) | (current_row >= 29);

  // assign vga_r = (lfsr[0] ^ lfsr[7]) & video_en;
  assign vga_r = color & video_en;
  // assign vga_g = (lfsr[1] ^ lfsr[12]) & video_en;
  // assign vga_b = (lfsr[2] ^ lfsr[5]) & video_en;
  // assign vga_g = mem_request & video_en;
  assign vga_g = 0 & video_en;
  //assign vga_b = (mem_request_complete | (pixel_x == 0) | (pixel_y == 0)) & video_en;
  // assign vga_b = ((pixel_x == 0) | (pixel_y == 0) & (current_col < 40)) & video_en;
  assign vga_b = 0 & video_en;

  assign vga_vs = scanline >= 2;
  assign vga_hs = (ctr < 2700) || (ctr > 3000);

  always @(posedge clk_100mhz) begin
    if (ena) begin
      if (!rst_n) begin
        ctr <= 0;
        scanline <= 0;
        line_flip <= 0;
        line_ctr <= 0;
        line_ptr <= 0;
        lfsr <= 1;
        video_mem_address <= 0;
      end else begin
        lfsr <= {lfsr[30:0], lfsr[31] ^ lfsr[21] ^ lfsr[1] ^ lfsr[0]};
        ctr <= ctr + 1;

        if (ctr >= 3200) begin
          ctr <= 0;
          scanline <= scanline < 524 ? scanline + 1 : 0;
          if (offset_scanline[3:0] == 4'b1111) begin
            line_flip <= !line_flip;
            line_ctr <= current_row;
            line_ptr <= 0;
          end
        end

        // Fetch the next line of characters.
        if ((line_ptr < 20) && (!video_mem_request) && (!video_mem_request_complete)) begin
          video_mem_address <= 40 * line_ctr + 2 * line_ptr;
          // video_mem_write_enable <= lfsr[0] & lfsr[1] & lfsr[2] & lfsr[3] & lfsr[4]; // FIXME: Do a random mixture of reads and writes.
          // video_mem_write_value <= lfsr[15:0];
          //video_mem_write_value <= video_mem_address;
          // video_mem_write_value <= 8'hc5;
          video_mem_write_enable <= 0;
          video_mem_request <= 1;
          line_ptr <= line_ptr + 1;
        end
        if (video_mem_request_complete) begin
          video_mem_request <= 0;
          if (line_flip) begin
            line_buffer1[line_ptr - 1] <= video_mem_read_value;
          end else begin
            line_buffer2[line_ptr - 1] <= video_mem_read_value;
          end
        end
      end
    end
  end
endmodule
