`define SRAM_ADDRESS_SIZE 17
`define SRAM_ADDRESS_IGNORED_BITS 7
`define MEMORY_WORD_SIZE 16

module memory_controller (
  input  wire                              ena,
  input  wire                              clk,
  input  wire                              rst_n,
  input  wire [`SRAM_ADDRESS_SIZE - 1 : 0] mem_address,
  input  wire [`MEMORY_WORD_SIZE - 1 : 0]  mem_write_value,
  input  wire                              mem_write_enable,
  output reg  [`MEMORY_WORD_SIZE - 1 : 0]  mem_read_value,
  input  wire                              mem_request,
  output reg                               mem_request_complete,
  output reg                               sram_cs_n,
  output reg                               sram_si,
  input  wire                              sram_so
);
  reg [11:0] counter;

  always @(posedge clk) begin
    if (ena) begin
      if (!rst_n) begin
        counter <= 0;
        sram_cs_n <= 1;
      end else begin
        if (mem_request) begin
          sram_cs_n <= 0;
          // The first seven bits are always 0, 0, 0, 0, 0, 0, 1
          if (counter < 6) begin
            sram_si <= 0;
          end else if (counter == 6) begin
            sram_si <= 1;
          end else if (counter == 7) begin
            // Then the eighth bit is 0 if we're writing, 1 if we're reading.
            sram_si <= !mem_write_enable;
          end else if (counter < 8 + `SRAM_ADDRESS_IGNORED_BITS) begin
            sram_si <= 0;
            // sram_si <= 1;
          end else if (counter < 32) begin
            // Then the next 17 bits are the address.
            //sram_si <= mem_address[`SRAM_ADDRESS_SIZE - (counter - 8 - `SRAM_ADDRESS_IGNORED_BITS) - 1];
            sram_si <= mem_address[counter - 8 - `SRAM_ADDRESS_IGNORED_BITS];
          end else if (counter < 32 + `MEMORY_WORD_SIZE) begin
            if (mem_write_enable) begin
              // Finally we send the bits to write, if relevant.
              sram_si <= mem_write_value[counter - 32];
            end else begin
              // Otherwise we read the bits.
              // $display("Reading bit %d = %d", counter - 32, sram_so);
              mem_read_value[counter - 32] <= sram_so;
            end
          end

          if (counter < 32 + `MEMORY_WORD_SIZE) begin
            counter <= counter + 1;
          end else begin
            counter <= 32 + `MEMORY_WORD_SIZE;
            mem_request_complete <= 1;
            sram_cs_n <= 1;
          end
        end else begin
          counter <= 0;
          mem_request_complete <= 0;
        end
      end
    end else begin
      sram_cs_n <= 1;
    end
  end
endmodule

module font_rom(
  input wire [7:0] char,
  input wire [3:0] pixel_x,
  input wire [3:0] pixel_y,
  output wire color
);
  assign color = char[{pixel_y[3], pixel_y[2], pixel_x[3]}];
  // reg [255:0] font [0:95];
  // initial begin
  //   font[0] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  //   font[1] = 256'b0000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000;
  //   font[2] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011000000000011001100000000001100110000000000110011000;
  //   font[3] = 256'b0000000000000000000000000000000000000001100110000000000110011000000000011001100000000001100110000000011111111110000001111111111000000001100110000000000110011000000001111111111000000111111111100000000110011000000000011001100000000001100110000000000110011000;
  //   font[4] = 256'b0000000000000000000000000000000000000000011000000000000001100000000000011111111000000011111111100000011001100000000001100110000000000011111111000000000111111110000000000110011000000000011001100000011111111110000001111111110000000000011000000000000001100000;
  //   font[5] = 256'b0000000000000000000000000000000000000111100001100000011110000110000001111000011000000111100011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100011110000001100001111000000110000111100000011000011110;
  //   font[6] = 256'b0000000000000000000000000000000000000010011111000000001111111110000000111100011000000011110001100000001111100110000000100111111000000000001111000000000000111100000000000111111000000000011001100000000001100110000000000110011000000000001111100000000000011100;
  //   font[7] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000000011000000000000001100000;
  //   font[8] = 256'b0000000000000000000000000000000000000001110000000000000111100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000001111000000000000111000000;
  //   font[9] = 256'b0000000000000000000000000000000000000000000110000000000000111000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000001110000000000000011000;
  //   font[10] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011000000000011001100000000000111100000000000011110000000001111111111000000111111111100000000011110000000000001111000000000001100110000000000110011000;
  //   font[11] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000011000000000000001100000000000000110000000000111111111100000011111111110000000000110000000000000011000000000000001100000000000000110000000000000000000000000000000000000;
  //   font[12] = 256'b0000000000011000000000000011100000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  //   font[13] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  //   font[14] = 256'b0000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  //   font[15] = 256'b0000000000000000000000000000000000000000000001100000000000000110000000000000011000000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000001100000000000000110000000000000011000000000;
  //   font[16] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000011110000001100011111000000110011101100000011011100110000001111100011000000111100001100000011100000110000001100000011000000011111111100000000111111100;
  //   font[17] = 256'b0000000000000000000000000000000000000001111110000000000111111000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001111000000000000111100000000000011100000000000001100000;
  //   font[18] = 256'b0000000000000000000000000000000000000111111111100000011111111110000000000001110000000000001110000000000001110000000000001110000000000001110000000000001110000000000001110000000000000110000000000000011000000110000001100000011000000011111111100000000111111100;
  //   font[19] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000000000001100000000000000011111000000000001111100000000001100000000000000110000000000000011000000110000001100000011000000011111111100000000111111100;
  //   font[20] = 256'b0000000000000000000000000000000000000001100000000000000110000000000000011000000000000001100000000000011111111110000001111111111000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100000000000000110000000;
  //   font[21] = 256'b0000000000000000000000000000000000000001111111100000001111111110000001100000000000000110000000000000011000000000000001100000000000000011111111100000000111111110000000000000011000000000000001100000000000000110000000000000011000000011111111100000001111111110;
  //   font[22] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111110000000000000011000000000000001100000000000000110000000000000011000000001111111100000000111111100;
  //   font[23] = 256'b0000000000000000000000000000000000000000000000100000000000000110000000000000110000000000000111000000000000111000000000000111000000000000111000000000000111000000000000111000000000000011000000000000001100000000000000110000000000000011111111100000001111111110;
  //   font[24] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000001111111100000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111100;
  //   font[25] = 256'b0000000000000000000000000000000000000001111111100000001111111110000001100000000000000110000000000000011000000000000001100000000000000111111111000000011111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111100;
  //   font[26] = 256'b0000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000011110000000000001111000000000000111100000000000000000000000000000000000;
  //   font[27] = 256'b0000000000011000000000000011100000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000011110000000000001111000000000000111100000000000000000000000000000000000;
  //   font[28] = 256'b0000000000000000000000000000000000000000100000000000000011000000000000000110000000000000001100000000000000111000000000000001110000000000000011100000000000001110000000000001110000000000001110000000000000110000000000000110000000000000110000000000000010000000;
  //   font[29] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000000000000000000000000000000000000001111111111000000111111111100000000000000000000000000000000000000000000000000000000000000000;
  //   font[30] = 256'b0000000000000000000000000000000000000000000110000000000000111000000000000111000000000000111000000000000111000000000000011000000000000011000000000000001100000000000000011000000000000001110000000000000011100000000000000111000000000000001110000000000000011000;
  //   font[31] = 256'b0000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000000001100000000000001110000000000001110000000000001110000000000001110000000000000110000000000000011000000110000001100000011000000011111111100000000111111100;
  //   font[32] = 256'b0000000000000000000000000000000000000111111111000000011111111110000000000000011000000000000001100000000111000110000000111110011000000110011001100000011001100110000001111110011000000111110001100000011000000110000001100000011000000011111111100000000111111100;
  //   font[33] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000111111111100000011111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111100;
  //   font[34] = 256'b0000000000000000000000000000000000000001111111100000001111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000001111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111110;
  //   font[35] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000011000000110000001100000011000000011111111100000000111111100;
  //   font[36] = 256'b0000000000000000000000000000000000000001111111100000001111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111110;
  //   font[37] = 256'b0000000000000000000000000000000000000011111111100000001111111110000000000000011000000000000001100000000000000110000000000000011000000000111111100000000011111110000000000000011000000000000001100000000000000110000000000000011000000011111111100000001111111110;
  //   font[38] = 256'b0000000000000000000000000000000000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000111111100000000011111110000000000000011000000000000001100000000000000110000000000000011000000011111111100000001111111110;
  //   font[39] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000110000001100000011000000111100001100000011110000110000000000000011000000000000001100000011000000110000001100000011000000011111111100000000111111100;
  //   font[40] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000111111111100000011111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110;
  //   font[41] = 256'b0000000000000000000000000000000000000001111110000000000111111000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000001111110000000000111111000;
  //   font[42] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000;
  //   font[43] = 256'b0000000000000000000000000000000000000010000001100000001100000110000000011000011000000001110001100000000011100110000000000111111000000000001111100000000000111110000000000111011000000000111001100000000011000110000000011000011000000011000001100000001000000110;
  //   font[44] = 256'b0000000000000000000000000000000000000011111111100000001111111110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110;
  //   font[45] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100110011000000110111101100000011111111110000001111001111000000111000011100000011000000110;
  //   font[46] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001110000011000000111100001100000011111000110000001101110011000000110011101100000011000111110000001100001111000000110000011100000011000000110;
  //   font[47] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111100;
  //   font[48] = 256'b0000000000000000000000000000000000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000001111111100000001111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111110;
  //   font[49] = 256'b0000000000000000000000000000000000000110011111000000011111111110000000111100011000000011110001100000011111100110000001100110011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111100;
  //   font[50] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000011111111100000001111111110000001100000011000000110000001100000011000000110000001100000011000000011111111100000000111111110;
  //   font[51] = 256'b0000000000000000000000000000000000000011111111000000001111111110000001100000011000000110000001100000011000000000000001100000000000000011111111000000000111111110000000000000011000000000000001100000011000000110000001100000011000000011111111100000000111111100;
  //   font[52] = 256'b0000000000000000000000000000000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000111111111100000011111111110;
  //   font[53] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110;
  //   font[54] = 256'b0000000000000000000000000000000000000000011000000000000011110000000000011111100000000011100111000000011100001110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110;
  //   font[55] = 256'b0000000000000000000000000000000000000001110111000000001111111110000001100110011000000110011001100000011001100110000001100110011000000110011001100000011001100110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110;
  //   font[56] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000111000011100000001110011100000000011111100000000000111100000000000011110000000000011111100000000011100111000000011100001110000001100000011000000110000001100000011000000110;
  //   font[57] = 256'b0000000000000000000000000000000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000011110000000000011111100000000011100111000000011100001110000001100000011000000110000001100000011000000110;
  //   font[58] = 256'b0000000000000000000000000000000000000011111111100000001111111110000000000000011000000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000011100000000000001100000000000000111111111000000011111111100;
  //   font[59] = 256'b0000000000000000000000000000000000000001111000000000000111100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000001111000000000000111100000;
  //   font[60] = 256'b0000000000000000000000000000000000000110000000000000011000000000000001100000000000000111000000000000001110000000000000011100000000000000111000000000000001110000000000000011100000000000000111000000000000001110000000000000011000000000000001100000000000000110;
  //   font[61] = 256'b0000000000000000000000000000000000000000011110000000000001111000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011110000000000001111000;
  //   font[62] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000111000011100000001110011100000000011111100000000000111100000000000001100000;
  //   font[63] = 256'b0000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  //   font[64] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000011100000000000000111000000000000001100000;
  //   font[65] = 256'b0000000000000000000000000000000000000111111111000000011111111110000001100000011000000110000001100000011111111110000001111111110000000110000000000000011000000000000000111111100000000001111110000000000000000000000000000000000000000000000000000000000000000000;
  //   font[66] = 256'b0000000000000000000000000000000000000001111111100000001111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000000111111111000000001111111100000000000000110000000000000011000000000000001100000000000000110;
  //   font[67] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000000000000110000000000000011000000110000001100000011000000110000000111111111000000001111111000000000000000000000000000000000000000000000000000000000000000000;
  //   font[68] = 256'b0000000000000000000000000000000000000111111111000000011111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001111111111000000111111111000000011000000000000001100000000000000110000000000000011000000000;
  //   font[69] = 256'b0000000000000000000000000000000000000001111111000000000111111110000000000000011000000000000001100000011111111110000001111111111000000110000001100000011000000110000000111111111000000001111111000000000000000000000000000000000000000000000000000000000000000000;
  //   font[70] = 256'b0000000000000000000000000000000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000011111100000000001111110000000000001100000000000000110000000000011111000000000001111000000;
  //   font[71] = 256'b0000000111111000000000111111100000000110000000000000011000000000000001111111110000000111111111100000011000000110000001100000011000000110000001100000011000000110000001111111111000000111111111000000000000000000000000000000000000000000000000000000000000000000;
  //   font[72] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000000111111111000000001111111100000000000000110000000000000011000000000000001100000000000000110;
  //   font[73] = 256'b0000000000000000000000000000000000000001111110000000000111111000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000111100000000000011110000000000000000000000000000000000000000000011000000000000001100000;
  //   font[74] = 256'b0000000001111100000000001111111000000001100001100000000110000110000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011110000000000001111000000000000000000000000000000000000000000001100000000000000110000000;
  //   font[75] = 256'b0000000000000000000000000000000000000010000110000000001100011000000000111001100000000001111110000000000011111000000000001111100000000001110110000000001110011000000000110001100000000010000110000000000000011000000000000001100000000000000110000000000000011000;
  //   font[76] = 256'b0000000000000000000000000000000000000001111110000000000111111000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011110000000000001111000;
  //   font[77] = 256'b0000000000000000000000000000000000000110011001100000011001100110000001100110011000000110011001100000011001100110000001100110011000000110011001100000011001100110000000111111111000000001100111100000000000000000000000000000000000000000000000000000000000000000;
  //   font[78] = 256'b0000000000000000000000000000000000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000000111111111000000001111111100000000000000000000000000000000000000000000000000000000000000000;
  //   font[79] = 256'b0000000000000000000000000000000000000001111111000000001111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000000111111111000000001111111000000000000000000000000000000000000000000000000000000000000000000;
  //   font[80] = 256'b0000000000000110000000000000011000000000000001100000000000000110000000011111111000000011111111100000011000000110000001100000011000000110000001100000011000000110000000111111111000000001111111100000000000000000000000000000000000000000000000000000000000000000;
  //   font[81] = 256'b0000011000000000000001100000000000000110000000000000011000000000000001111111110000000111111111100000011000000110000001100000011000000110000001100000011000000110000001111111111000000111111111000000000000000000000000000000000000000000000000000000000000000000;
  //   font[82] = 256'b0000000000000000000000000000000000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000110000110000000011000011000000000111111100000000001111110000000000000000000000000000000000000000000000000000000000000000000;
  //   font[83] = 256'b0000000000000000000000000000000000000001111111100000001111111110000001100000000000000110000000000000001111111100000000011111111000000000000001100000000000000110000001111111111000000111111111000000000000000000000000000000000000000000000000000000000000000000;
  //   font[84] = 256'b0000000000000000000000000000000000000111110000000000011111100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000001111111100000000111111110000000000001100000000000000110000000000000011000000000000001100000;
  //   font[85] = 256'b0000000000000000000000000000000000000111111111000000011111111110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000000000000000000000000000000000000000000000000000000000000000;
  //   font[86] = 256'b0000000000000000000000000000000000000000011000000000000011110000000000011111100000000011100111000000011100001110000001100000011000000110000001100000011000000110000001100000011000000110000001100000000000000000000000000000000000000000000000000000000000000000;
  //   font[87] = 256'b0000000000000000000000000000000000000001110111000000001111111110000001100110011000000110011001100000011001100110000001100110011000000110011001100000011001100110000001100000011000000110000001100000000000000000000000000000000000000000000000000000000000000000;
  //   font[88] = 256'b0000000000000000000000000000000000000110000001100000011100001110000000111001110000000001111110000000000011110000000000001111000000000001111110000000001110011100000001110000111000000110000001100000000000000000000000000000000000000000000000000000000000000000;
  //   font[89] = 256'b0000000111111000000000111111100000000110000000000000011000000000000001111111110000000111111111100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000000000000000000000000000000000000000000000000000000000000000;
  //   font[90] = 256'b0000000000000000000000000000000000000111111111100000011111111110000000000001110000000000001110000000000001110000000000001110000000000001110000000000001110000000000001111111111000000111111111100000000000000000000000000000000000000000000000000000000000000000;
  //   font[91] = 256'b0000000000000000000000000000000000000001110000000000000111100000000000000110000000000000011000000000000001100000000000000110000000000000001110000000000000111000000000000110000000000000011000000000000001100000000000000110000000000001111000000000000111000000;
  //   font[92] = 256'b0000000000000000000000000000000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000;
  //   font[93] = 256'b0000000000000000000000000000000000000000000110000000000000111000000000000110000000000000011000000000000001100000000000000110000000000001110000000000000111100000000000000110000000000000011000000000000001100000000000000110000000000000001110000000000000011000;
  //   font[94] = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000011111000000000011001100110000001100110011000000000001111000000000000011100;
  //   font[95] = 256'b0000000000000000000000000000000000000111111111100000011111111110000001111111111000000111111111100000011111111110000001111111111000000111111111100000011111111110000001111111111000000111111111100000011111111110000001111111111000000111111111100000011111111110;
  // end
  // assign color = ((char >= 32) && (char < 96)) ? font[char - 32][pixel_y * 16 + pixel_x] : pixel_x ^ pixel_y;
endmodule

// PMOD0 is the output for the VGA.
// PMOD1 is the input/output for the SRAM.
//   PMOD1[0]: ~CS
//   PMOD1[1]: SO
//   PMOD1[2]: SIO2
//   PMOD1[3]: SI
//   PMOD1[4]: SCK
//   PMOD1[5]: ~HOLD/SIO3

module micro1 (
  input  wire [7:0] ui_in,      // dedicated inputs
  output wire [7:0] uo_out,     // dedicated outputs
  input  wire [7:0] uio_in,     // bidirectional input path
  output wire [7:0] uio_out,    // bidirectional output path
  output wire [7:0] uio_oe,     // bidir output enable (high=out)
  input  wire       ena,        // high when enabled
  input  wire       clk_100mhz, // clock
  input  wire       rst_n       // reset negated (low to reset)
);
  wire vga_r = uo_out[0];
  wire vga_g = uo_out[1];
  wire vga_b = uo_out[2];
  wire vga_hs = uo_out[3];
  wire vga_vs = uo_out[4];

  reg [`SRAM_ADDRESS_SIZE - 1 : 0] mem_address;
  reg [`MEMORY_WORD_SIZE - 1 : 0]  mem_write_value;
  reg                              mem_write_enable;
  reg [`MEMORY_WORD_SIZE - 1 : 0]  mem_read_value;
  reg                              mem_request;
  reg                              mem_request_complete;

  // Set output directions.
  assign uio_oe[0] = 1;
  assign uio_oe[1] = 0;
  assign uio_oe[2] = 1; // We're pulling up, so output.
  assign uio_oe[3] = 1;
  assign uio_oe[4] = 1;
  assign uio_oe[5] = 1; // We're pulling up, so output.
  // Assign pull-up values.
  assign uio_out[2] = 1;
  assign uio_out[5] = 1;

  reg [3:0] mem_controller_clock_divider = 0;
  always @(posedge clk_100mhz) begin
    mem_controller_clock_divider <= mem_controller_clock_divider + 1;
  end

  // Assign the serial clock.
  assign uio_out[4] = !(mem_controller_clock_divider[3] ^ mem_controller_clock_divider[2]);

  memory_controller memory_controller_inst(
    .ena(ena),
    .clk(mem_controller_clock_divider[3]),
    .rst_n(rst_n),
    .mem_address(mem_address),
    .mem_write_value(mem_write_value),
    .mem_write_enable(mem_write_enable),
    .mem_read_value(mem_read_value),
    .mem_request(mem_request),
    .mem_request_complete(mem_request_complete),
    .sram_cs_n(uio_out[0]),
    .sram_si(uio_out[3]),
    .sram_so(uio_in[1])
  );

  reg [23:0] ctr = 0;
  reg [15:0] scanline = 0;
  reg [31:0] lfsr = 1;

  reg [15:0] line_buffer1 [0:19];
  reg [15:0] line_buffer2 [0:19];
  reg line_flip = 0;
  reg [5:0] line_ctr = 0;
  reg [4:0] line_ptr = 0;

  reg mem_fill = 0;

  wire video_en = (scanline >= 35) && (scanline < 515) && (ctr < 2700);

  // We now figure out which character we're at.
  wire [9:0] offset_scanline = scanline - 35;
  wire [4:0] current_row = offset_scanline[8:4];
  wire [3:0] pixel_y = offset_scanline[3:0];
  // Each pixel is 4 cycles long.
  wire [6:0] current_col = ctr[12:6];
  wire [3:0] pixel_x = ctr[5:2];

  wire [15:0] current_char_pair = current_col >= 40 ? 0 : (line_flip ? line_buffer2[current_col >> 1] : line_buffer1[current_col >> 1]);
  wire [7:0] current_char = current_col[0] ? current_char_pair[7:0] : current_char_pair[15:8];

  wire color;
  font_rom font_rom_inst(
    .char(current_char),
    .pixel_x(pixel_x),
    .pixel_y(pixel_y),
    .color(color)
  );

  // We now interpret the character as a little 2x4 grid.
  // wire color = current_char[{pixel_y[3], pixel_y[2], pixel_x[3]}];
  //wire color = (current_col >= 39) | (current_row >= 29);

  // assign vga_r = (lfsr[0] ^ lfsr[7]) & video_en;
  assign vga_r = color & video_en;
  // assign vga_g = (lfsr[1] ^ lfsr[12]) & video_en;
  // assign vga_b = (lfsr[2] ^ lfsr[5]) & video_en;
  // assign vga_g = mem_request & video_en;
  assign vga_g = 0 & video_en;
  //assign vga_b = (mem_request_complete | (pixel_x == 0) | (pixel_y == 0)) & video_en;
  // assign vga_b = ((pixel_x == 0) | (pixel_y == 0) & (current_col < 40)) & video_en;
  assign vga_b = 0 & video_en;

  assign vga_vs = scanline >= 2;
  assign vga_hs = (ctr < 2700) || (ctr > 3000);

  always @(posedge clk_100mhz) begin
    if (ena) begin
      if (!rst_n) begin
        ctr <= 0;
        scanline <= 0;
        line_flip <= 0;
        line_ctr <= 0;
        line_ptr <= 0;
        lfsr <= 1;
        mem_fill <= 1;
        mem_address <= 0;
      end else begin
        lfsr <= {lfsr[30:0], lfsr[31] ^ lfsr[21] ^ lfsr[1] ^ lfsr[0]};
        ctr <= ctr + 1;

        if (ctr >= 3200) begin
          ctr <= 0;
          scanline <= scanline < 524 ? scanline + 1 : 0;
          if (offset_scanline[3:0] == 4'b1111) begin
            line_flip <= !line_flip;
            line_ctr <= current_row;
            line_ptr <= 0;
          end
        end

        if (mem_fill) begin
          // Begin filling memory with characters.
          if (!mem_request) begin
            mem_address <= mem_address + 1;
            mem_write_value <= lfsr[15:0];
            mem_write_enable <= 1;
            mem_request <= 1;
          end
          if (mem_request_complete) begin
            mem_request <= 0;
            if (mem_address >= 1200) begin
              mem_fill <= 0;
            end
          end
        end else begin
          // Otherwise, fetch the next line of characters.
          if ((line_ptr < 20) && (!mem_request) && (!mem_request_complete)) begin
            mem_address <= 40 * line_ctr + 2 * line_ptr;
            mem_write_enable <= lfsr[0] & lfsr[1] & lfsr[2] & lfsr[3] & lfsr[4]; // FIXME: Do a random mixture of reads and writes.
            mem_write_value <= lfsr[15:0];
            //mem_write_value <= mem_address;
            // mem_write_value <= 8'hc5;
            // mem_write_enable <= 0;
            mem_request <= 1;
            line_ptr <= line_ptr + 1;
          end
          if (mem_request_complete) begin
            mem_request <= 0;
            if (line_flip) begin
              line_buffer1[line_ptr - 1] <= mem_read_value;
            end else begin
              line_buffer2[line_ptr - 1] <= mem_read_value;
            end
          end

        end
      end
    end
  end
endmodule
